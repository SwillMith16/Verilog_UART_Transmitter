library verilog;
use verilog.vl_types.all;
entity tx_7seg_decoder_vlg_vec_tst is
end tx_7seg_decoder_vlg_vec_tst;
