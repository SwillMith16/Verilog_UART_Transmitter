library verilog;
use verilog.vl_types.all;
entity tx_bit_counter_vlg_vec_tst is
end tx_bit_counter_vlg_vec_tst;
