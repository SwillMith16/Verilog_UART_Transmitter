library verilog;
use verilog.vl_types.all;
entity tx_3to4_bus_expansion_vlg_vec_tst is
end tx_3to4_bus_expansion_vlg_vec_tst;
